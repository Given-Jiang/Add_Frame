-- Add_Frame_GN_Add_Frame_Add_Frame_Module_CTRL_DECODER.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.25.10:37:28

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Add_Frame_GN_Add_Frame_Add_Frame_Module_CTRL_DECODER is
	port (
		decoder_col : out std_logic_vector(15 downto 0);                    -- decoder_col.wire
		decoder_row : out std_logic_vector(15 downto 0);                    -- decoder_row.wire
		height      : out std_logic_vector(15 downto 0);                    --      height.wire
		data        : in  std_logic_vector(23 downto 0) := (others => '0'); --        data.wire
		sop         : in  std_logic                     := '0';             --         sop.wire
		width       : out std_logic_vector(15 downto 0);                    --       width.wire
		Clock       : in  std_logic                     := '0';             --       Clock.clk
		aclr        : in  std_logic                     := '0'              --            .reset
	);
end entity Add_Frame_GN_Add_Frame_Add_Frame_Module_CTRL_DECODER;

architecture rtl of Add_Frame_GN_Add_Frame_Add_Frame_Module_CTRL_DECODER is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_cast_GNED3D3FSF is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNED3D3FSF;

	component alt_dspbuilder_cast_GNYDD6MCZ4 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNYDD6MCZ4;

	component alt_dspbuilder_cast_GNHBD5Z3AF is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNHBD5Z3AF;

	component alt_dspbuilder_cast_GN76IOUHQH is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GN76IOUHQH;

	component alt_dspbuilder_cast_GNMU5M7DX7 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNMU5M7DX7;

	component alt_dspbuilder_cast_GNI42JW6WW is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNI42JW6WW;

	component alt_dspbuilder_bus_concat_GNAUBM7IRL is
		generic (
			widthB : natural := 8;
			widthA : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNAUBM7IRL;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_bus_concat_GNBH75ZTOD is
		generic (
			widthB : natural := 8;
			widthA : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNBH75ZTOD;

	component alt_dspbuilder_bus_concat_GNXPBV3I7L is
		generic (
			widthB : natural := 8;
			widthA : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNXPBV3I7L;

	component alt_dspbuilder_port_GNBO6OMO5Y is
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNBO6OMO5Y;

	component alt_dspbuilder_if_statement_GNURIZNNI4 is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                       -- wire
			a    : in  std_logic_vector(2 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(2 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNURIZNNI4;

	component alt_dspbuilder_constant_GNP7P5YZV2 is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(2 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNP7P5YZV2;

	component alt_dspbuilder_logical_bit_op_GNKUBZL4TE is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNKUBZL4TE;

	component alt_dspbuilder_logical_bit_op_GNUQ2R64DV is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNUQ2R64DV;

	component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V;

	component alt_dspbuilder_delay_GNVCBR7UZP is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNVCBR7UZP;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_counter_GNW5IG44CT is
		generic (
			use_usr_aclr : string  := "false";
			use_ena      : string  := "false";
			use_cin      : string  := "false";
			use_sset     : string  := "false";
			ndirection   : natural := 1;
			svalue       : string  := "0";
			use_sload    : string  := "false";
			use_sclr     : string  := "false";
			use_cout     : string  := "false";
			modulus      : integer := 256;
			use_cnt_ena  : string  := "false";
			width        : natural := 8;
			use_aset     : string  := "false";
			use_aload    : string  := "false";
			avalue       : string  := "0"
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			aload     : in  std_logic                          := 'X';             -- wire
			aset      : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cnt_ena   : in  std_logic                          := 'X';             -- wire
			cout      : out std_logic;                                             -- wire
			data      : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			direction : in  std_logic                          := 'X';             -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			q         : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr      : in  std_logic                          := 'X';             -- wire
			sload     : in  std_logic                          := 'X';             -- wire
			sset      : in  std_logic                          := 'X';             -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_counter_GNW5IG44CT;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_delay_GNGQ56ZS4N is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNGQ56ZS4N;

	component alt_dspbuilder_decoder_GNSCEXJCJK is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNSCEXJCJK;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_cast_GNSB3OXIQS is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			output : out std_logic                                        -- wire
		);
	end component alt_dspbuilder_cast_GNSB3OXIQS;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	signal delay5sclrgnd_output_wire         : std_logic;                     -- Delay5sclrGND:output -> Delay5:sclr
	signal delay4sclrgnd_output_wire         : std_logic;                     -- Delay4sclrGND:output -> Delay4:sclr
	signal delay3sclrgnd_output_wire         : std_logic;                     -- Delay3sclrGND:output -> Delay3:sclr
	signal delay1sclrgnd_output_wire         : std_logic;                     -- Delay1sclrGND:output -> Delay1:sclr
	signal decodersclrgnd_output_wire        : std_logic;                     -- DecodersclrGND:output -> Decoder:sclr
	signal decoderenavcc_output_wire         : std_logic;                     -- DecoderenaVCC:output -> Decoder:ena
	signal bus_concatenation3_output_wire    : std_logic_vector(7 downto 0);  -- Bus_Concatenation3:output -> Bus_Concatenation4:a
	signal bus_concatenation5_output_wire    : std_logic_vector(7 downto 0);  -- Bus_Concatenation5:output -> Bus_Concatenation1:a
	signal bus_concatenation4_output_wire    : std_logic_vector(11 downto 0); -- Bus_Concatenation4:output -> Bus_Concatenation6:a
	signal bus_concatenation7_output_wire    : std_logic_vector(7 downto 0);  -- Bus_Concatenation7:output -> Bus_Concatenation8:a
	signal bus_concatenation8_output_wire    : std_logic_vector(11 downto 0); -- Bus_Concatenation8:output -> Bus_Concatenation9:a
	signal data_0_output_wire                : std_logic_vector(23 downto 0); -- data_0:output -> [Bus_Conversion1:input, Bus_Conversion2:input, Bus_Conversion3:input, Decoder:data]
	signal bus_conversion1_output_wire       : std_logic_vector(3 downto 0);  -- Bus_Conversion1:output -> Bus_Concatenation5:b
	signal bus_conversion10_output_wire      : std_logic_vector(3 downto 0);  -- Bus_Conversion10:output -> Bus_Concatenation8:b
	signal bus_conversion11_output_wire      : std_logic_vector(3 downto 0);  -- Bus_Conversion11:output -> Bus_Concatenation9:b
	signal bus_conversion2_output_wire       : std_logic_vector(3 downto 0);  -- Bus_Conversion2:output -> Bus_Concatenation5:a
	signal bus_conversion3_output_wire       : std_logic_vector(3 downto 0);  -- Bus_Conversion3:output -> Bus_Concatenation1:b
	signal bus_conversion4_output_wire       : std_logic_vector(3 downto 0);  -- Bus_Conversion4:output -> Bus_Concatenation3:a
	signal bus_conversion5_output_wire       : std_logic_vector(3 downto 0);  -- Bus_Conversion5:output -> Bus_Concatenation3:b
	signal bus_conversion6_output_wire       : std_logic_vector(3 downto 0);  -- Bus_Conversion6:output -> Bus_Concatenation4:b
	signal bus_conversion7_output_wire       : std_logic_vector(3 downto 0);  -- Bus_Conversion7:output -> Bus_Concatenation6:b
	signal bus_conversion8_output_wire       : std_logic_vector(3 downto 0);  -- Bus_Conversion8:output -> Bus_Concatenation7:a
	signal bus_conversion9_output_wire       : std_logic_vector(3 downto 0);  -- Bus_Conversion9:output -> Bus_Concatenation7:b
	signal delay3_output_wire                : std_logic_vector(11 downto 0); -- Delay3:output -> [Bus_Conversion4:input, Bus_Conversion5:input, Bus_Conversion6:input]
	signal delay4_output_wire                : std_logic_vector(11 downto 0); -- Delay4:output -> [Bus_Conversion7:input, Bus_Conversion8:input, Bus_Conversion9:input, Delay3:input]
	signal bus_concatenation1_output_wire    : std_logic_vector(11 downto 0); -- Bus_Concatenation1:output -> Delay5:input
	signal delay5_output_wire                : std_logic_vector(11 downto 0); -- Delay5:output -> [Bus_Conversion10:input, Bus_Conversion11:input, Bus_Conversion12:input, Delay4:input]
	signal constant2_output_wire             : std_logic_vector(2 downto 0);  -- Constant2:output -> If_Statement:a
	signal counter_q_wire                    : std_logic_vector(2 downto 0);  -- Counter:q -> If_Statement:b
	signal decoder_dec_wire                  : std_logic;                     -- Decoder:dec -> Logical_Bit_Operator:data0
	signal sop_0_output_wire                 : std_logic;                     -- sop_0:output -> Logical_Bit_Operator:data1
	signal logical_bit_operator_result_wire  : std_logic;                     -- Logical_Bit_Operator:result -> [Logical_Bit_Operator1:data0, cast221:input]
	signal if_statement_true_wire            : std_logic;                     -- If_Statement:true -> Logical_Bit_Operator1:data1
	signal logical_bit_operator1_result_wire : std_logic;                     -- Logical_Bit_Operator1:result -> Delay1:ena
	signal logical_bit_operator3_result_wire : std_logic;                     -- Logical_Bit_Operator3:result -> Counter:sclr
	signal bus_concatenation6_output_wire    : std_logic_vector(15 downto 0); -- Bus_Concatenation6:output -> [decoder_col_0:input, width_0:input]
	signal bus_concatenation9_output_wire    : std_logic_vector(15 downto 0); -- Bus_Concatenation9:output -> [decoder_row_0:input, height_0:input]
	signal delay1_output_wire                : std_logic_vector(0 downto 0);  -- Delay1:output -> [cast217:input, cast218:input, cast219:input, cast220:input, cast222:input]
	signal cast217_output_wire               : std_logic;                     -- cast217:output -> Counter:cnt_ena
	signal cast218_output_wire               : std_logic;                     -- cast218:output -> Delay3:ena
	signal cast219_output_wire               : std_logic;                     -- cast219:output -> Delay4:ena
	signal cast220_output_wire               : std_logic;                     -- cast220:output -> Delay5:ena
	signal cast221_output_wire               : std_logic_vector(0 downto 0);  -- cast221:output -> Delay1:input
	signal cast222_output_wire               : std_logic;                     -- cast222:output -> Logical_Bit_Operator3:data0
	signal clock_0_clock_output_reset        : std_logic;                     -- Clock_0:aclr_out -> [Bus_Concatenation1:aclr, Bus_Concatenation3:aclr, Bus_Concatenation4:aclr, Bus_Concatenation5:aclr, Bus_Concatenation6:aclr, Bus_Concatenation7:aclr, Bus_Concatenation8:aclr, Bus_Concatenation9:aclr, Counter:aclr, Decoder:aclr, Delay1:aclr, Delay3:aclr, Delay4:aclr, Delay5:aclr]
	signal clock_0_clock_output_clk          : std_logic;                     -- Clock_0:clock_out -> [Bus_Concatenation1:clock, Bus_Concatenation3:clock, Bus_Concatenation4:clock, Bus_Concatenation5:clock, Bus_Concatenation6:clock, Bus_Concatenation7:clock, Bus_Concatenation8:clock, Bus_Concatenation9:clock, Counter:clock, Decoder:clock, Delay1:clock, Delay3:clock, Delay4:clock, Delay5:clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	bus_conversion1 : component alt_dspbuilder_cast_GNED3D3FSF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_0_output_wire,          --  input.wire
			output => bus_conversion1_output_wire  -- output.wire
		);

	bus_conversion12 : component alt_dspbuilder_cast_GNYDD6MCZ4
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay5_output_wire, --  input.wire
			output => open                -- output.wire
		);

	bus_conversion2 : component alt_dspbuilder_cast_GNHBD5Z3AF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_0_output_wire,          --  input.wire
			output => bus_conversion2_output_wire  -- output.wire
		);

	bus_conversion10 : component alt_dspbuilder_cast_GN76IOUHQH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay5_output_wire,           --  input.wire
			output => bus_conversion10_output_wire  -- output.wire
		);

	bus_conversion3 : component alt_dspbuilder_cast_GNMU5M7DX7
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_0_output_wire,          --  input.wire
			output => bus_conversion3_output_wire  -- output.wire
		);

	bus_conversion11 : component alt_dspbuilder_cast_GNI42JW6WW
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay5_output_wire,           --  input.wire
			output => bus_conversion11_output_wire  -- output.wire
		);

	bus_conversion4 : component alt_dspbuilder_cast_GN76IOUHQH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay3_output_wire,          --  input.wire
			output => bus_conversion4_output_wire  -- output.wire
		);

	bus_concatenation7 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => bus_conversion8_output_wire,    --          a.wire
			b      => bus_conversion9_output_wire,    --          b.wire
			output => bus_concatenation7_output_wire  --     output.wire
		);

	data_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => data,               --  input.wire
			output => data_0_output_wire  -- output.wire
		);

	bus_concatenation8 : component alt_dspbuilder_bus_concat_GNBH75ZTOD
		generic map (
			widthB => 4,
			widthA => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => bus_concatenation7_output_wire, --          a.wire
			b      => bus_conversion10_output_wire,   --          b.wire
			output => bus_concatenation8_output_wire  --     output.wire
		);

	bus_concatenation5 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => bus_conversion2_output_wire,    --          a.wire
			b      => bus_conversion1_output_wire,    --          b.wire
			output => bus_concatenation5_output_wire  --     output.wire
		);

	bus_concatenation6 : component alt_dspbuilder_bus_concat_GNXPBV3I7L
		generic map (
			widthB => 4,
			widthA => 12
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => bus_concatenation4_output_wire, --          a.wire
			b      => bus_conversion7_output_wire,    --          b.wire
			output => bus_concatenation6_output_wire  --     output.wire
		);

	bus_concatenation3 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => bus_conversion4_output_wire,    --          a.wire
			b      => bus_conversion5_output_wire,    --          b.wire
			output => bus_concatenation3_output_wire  --     output.wire
		);

	bus_concatenation4 : component alt_dspbuilder_bus_concat_GNBH75ZTOD
		generic map (
			widthB => 4,
			widthA => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => bus_concatenation3_output_wire, --          a.wire
			b      => bus_conversion6_output_wire,    --          b.wire
			output => bus_concatenation4_output_wire  --     output.wire
		);

	bus_concatenation1 : component alt_dspbuilder_bus_concat_GNBH75ZTOD
		generic map (
			widthB => 4,
			widthA => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => bus_concatenation5_output_wire, --          a.wire
			b      => bus_conversion3_output_wire,    --          b.wire
			output => bus_concatenation1_output_wire  --     output.wire
		);

	height_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => bus_concatenation9_output_wire, --  input.wire
			output => height                          -- output.wire
		);

	if_statement : component alt_dspbuilder_if_statement_GNURIZNNI4
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "(a<b)",
			number_inputs   => 2,
			width           => 3
		)
		port map (
			true => if_statement_true_wire, -- true.wire
			a    => constant2_output_wire,  --    a.wire
			b    => counter_q_wire          --    b.wire
		);

	constant2 : component alt_dspbuilder_constant_GNP7P5YZV2
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "001",
			width      => 3
		)
		port map (
			output => constant2_output_wire  -- output.wire
		);

	logical_bit_operator3 : component alt_dspbuilder_logical_bit_op_GNKUBZL4TE
		generic map (
			LogicalOp     => "AltNOT",
			number_inputs => 1
		)
		port map (
			result => logical_bit_operator3_result_wire, -- result.wire
			data0  => cast222_output_wire                --  data0.wire
		);

	logical_bit_operator1 : component alt_dspbuilder_logical_bit_op_GNUQ2R64DV
		generic map (
			LogicalOp     => "AltOR",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator1_result_wire, -- result.wire
			data0  => logical_bit_operator_result_wire,  --  data0.wire
			data1  => if_statement_true_wire             --  data1.wire
		);

	decoder_row_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => bus_concatenation9_output_wire, --  input.wire
			output => decoder_row                     -- output.wire
		);

	logical_bit_operator : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator_result_wire, -- result.wire
			data0  => decoder_dec_wire,                 --  data0.wire
			data1  => sop_0_output_wire                 --  data1.wire
		);

	width_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => bus_concatenation6_output_wire, --  input.wire
			output => width                           -- output.wire
		);

	decoder_col_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => bus_concatenation6_output_wire, --  input.wire
			output => decoder_col                     -- output.wire
		);

	delay5 : component alt_dspbuilder_delay_GNVCBR7UZP
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "000000000001",
			width      => 12
		)
		port map (
			input  => bus_concatenation1_output_wire, --      input.wire
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			output => delay5_output_wire,             --     output.wire
			sclr   => delay5sclrgnd_output_wire,      --       sclr.wire
			ena    => cast220_output_wire             --        ena.wire
		);

	delay5sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay5sclrgnd_output_wire  -- output.wire
		);

	counter : component alt_dspbuilder_counter_GNW5IG44CT
		generic map (
			use_usr_aclr => "false",
			use_ena      => "false",
			use_cin      => "false",
			use_sset     => "false",
			ndirection   => 1,
			svalue       => "1",
			use_sload    => "false",
			use_sclr     => "true",
			use_cout     => "false",
			modulus      => -1,
			use_cnt_ena  => "true",
			width        => 3,
			use_aset     => "false",
			use_aload    => "false",
			avalue       => "0"
		)
		port map (
			clock   => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr    => clock_0_clock_output_reset,        --           .reset
			cnt_ena => cast217_output_wire,               --    cnt_ena.wire
			sclr    => logical_bit_operator3_result_wire, --       sclr.wire
			q       => counter_q_wire,                    --          q.wire
			cout    => open                               --       cout.wire
		);

	delay4 : component alt_dspbuilder_delay_GNVCBR7UZP
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "000000000001",
			width      => 12
		)
		port map (
			input  => delay5_output_wire,         --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay4_output_wire,         --     output.wire
			sclr   => delay4sclrgnd_output_wire,  --       sclr.wire
			ena    => cast219_output_wire         --        ena.wire
		);

	delay4sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay4sclrgnd_output_wire  -- output.wire
		);

	delay3 : component alt_dspbuilder_delay_GNVCBR7UZP
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "000000000001",
			width      => 12
		)
		port map (
			input  => delay4_output_wire,         --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay3_output_wire,         --     output.wire
			sclr   => delay3sclrgnd_output_wire,  --       sclr.wire
			ena    => cast218_output_wire         --        ena.wire
		);

	delay3sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay3sclrgnd_output_wire  -- output.wire
		);

	sop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sop,               --  input.wire
			output => sop_0_output_wire  -- output.wire
		);

	bus_concatenation9 : component alt_dspbuilder_bus_concat_GNXPBV3I7L
		generic map (
			widthB => 4,
			widthA => 12
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => bus_concatenation8_output_wire, --          a.wire
			b      => bus_conversion11_output_wire,   --          b.wire
			output => bus_concatenation9_output_wire  --     output.wire
		);

	delay1 : component alt_dspbuilder_delay_GNGQ56ZS4N
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "1",
			width      => 1
		)
		port map (
			input  => cast221_output_wire,               --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay1_output_wire,                --     output.wire
			sclr   => delay1sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator1_result_wire  --        ena.wire
		);

	delay1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay1sclrgnd_output_wire  -- output.wire
		);

	bus_conversion9 : component alt_dspbuilder_cast_GNYDD6MCZ4
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay4_output_wire,          --  input.wire
			output => bus_conversion9_output_wire  -- output.wire
		);

	bus_conversion8 : component alt_dspbuilder_cast_GNI42JW6WW
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay4_output_wire,          --  input.wire
			output => bus_conversion8_output_wire  -- output.wire
		);

	decoder : component alt_dspbuilder_decoder_GNSCEXJCJK
		generic map (
			decode   => "000000000000000000001111",
			pipeline => 0,
			width    => 24
		)
		port map (
			clock => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset, --           .reset
			data  => data_0_output_wire,         --       data.wire
			dec   => decoder_dec_wire,           --        dec.wire
			sclr  => decodersclrgnd_output_wire, --       sclr.wire
			ena   => decoderenavcc_output_wire   --        ena.wire
		);

	decodersclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decodersclrgnd_output_wire  -- output.wire
		);

	decoderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoderenavcc_output_wire  -- output.wire
		);

	bus_conversion7 : component alt_dspbuilder_cast_GN76IOUHQH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay4_output_wire,          --  input.wire
			output => bus_conversion7_output_wire  -- output.wire
		);

	bus_conversion6 : component alt_dspbuilder_cast_GNYDD6MCZ4
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay3_output_wire,          --  input.wire
			output => bus_conversion6_output_wire  -- output.wire
		);

	bus_conversion5 : component alt_dspbuilder_cast_GNI42JW6WW
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay3_output_wire,          --  input.wire
			output => bus_conversion5_output_wire  -- output.wire
		);

	cast217 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire,  --  input.wire
			output => cast217_output_wire  -- output.wire
		);

	cast218 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire,  --  input.wire
			output => cast218_output_wire  -- output.wire
		);

	cast219 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire,  --  input.wire
			output => cast219_output_wire  -- output.wire
		);

	cast220 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire,  --  input.wire
			output => cast220_output_wire  -- output.wire
		);

	cast221 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator_result_wire, --  input.wire
			output => cast221_output_wire               -- output.wire
		);

	cast222 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire,  --  input.wire
			output => cast222_output_wire  -- output.wire
		);

end architecture rtl; -- of Add_Frame_GN_Add_Frame_Add_Frame_Module_CTRL_DECODER
