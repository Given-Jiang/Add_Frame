-- Add_Frame_GN.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.25.10:37:27

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Add_Frame_GN is
	port (
		Avalon_ST_Sink_data                                 : in  std_logic_vector(23 downto 0) := (others => '0'); --                                 Avalon_ST_Sink_data.wire
		Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_col : out std_logic_vector(15 downto 0);                    -- Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_col.wire
		Avalon_ST_Source_ready                              : in  std_logic                     := '0';             --                              Avalon_ST_Source_ready.wire
		Avalon_ST_Sink_valid                                : in  std_logic                     := '0';             --                                Avalon_ST_Sink_valid.wire
		Avalon_MM_Slave_writedata                           : in  std_logic_vector(31 downto 0) := (others => '0'); --                           Avalon_MM_Slave_writedata.wire
		Add_Frame_Add_Frame_Module_state                    : out std_logic_vector(2 downto 0);                     --                    Add_Frame_Add_Frame_Module_state.wire
		Avalon_ST_Sink_endofpacket                          : in  std_logic                     := '0';             --                          Avalon_ST_Sink_endofpacket.wire
		Avalon_ST_Source_valid                              : out std_logic;                                        --                              Avalon_ST_Source_valid.wire
		Clock                                               : in  std_logic                     := '0';             --                                               Clock.clk
		aclr                                                : in  std_logic                     := '0';             --                                                    .reset
		Add_Frame_Add_Frame_Module_row_counter              : out std_logic_vector(15 downto 0);                    --              Add_Frame_Add_Frame_Module_row_counter.wire
		Avalon_MM_Slave_address                             : in  std_logic_vector(2 downto 0)  := (others => '0'); --                             Avalon_MM_Slave_address.wire
		Avalon_MM_Slave_write                               : in  std_logic                     := '0';             --                               Avalon_MM_Slave_write.wire
		Avalon_ST_Sink_ready                                : out std_logic;                                        --                                Avalon_ST_Sink_ready.wire
		Avalon_ST_Sink_startofpacket                        : in  std_logic                     := '0';             --                        Avalon_ST_Sink_startofpacket.wire
		Add_Frame_Add_Frame_Module_frame_in                 : out std_logic_vector(0 downto 0);                     --                 Add_Frame_Add_Frame_Module_frame_in.wire
		Avalon_ST_Source_startofpacket                      : out std_logic;                                        --                      Avalon_ST_Source_startofpacket.wire
		Add_Frame_Add_Frame_Module_col_counter              : out std_logic_vector(15 downto 0);                    --              Add_Frame_Add_Frame_Module_col_counter.wire
		Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_row : out std_logic_vector(15 downto 0);                    -- Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_row.wire
		Avalon_ST_Source_endofpacket                        : out std_logic;                                        --                        Avalon_ST_Source_endofpacket.wire
		Avalon_ST_Source_data                               : out std_logic_vector(23 downto 0)                     --                               Avalon_ST_Source_data.wire
	);
end entity Add_Frame_GN;

architecture rtl of Add_Frame_GN is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_port_GNS2GDLO5E is
		port (
			input  : in  std_logic_vector(2 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(2 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNS2GDLO5E;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component Add_Frame_GN_Add_Frame_Add_Frame_Module is
		port (
			state                                               : out std_logic_vector(2 downto 0);                     -- wire
			writedata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_col : out std_logic_vector(15 downto 0);                    -- wire
			addr                                                : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- wire
			data_in                                             : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			data_out                                            : out std_logic_vector(23 downto 0);                    -- wire
			Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_row : out std_logic_vector(15 downto 0);                    -- wire
			col_counter                                         : out std_logic_vector(15 downto 0);                    -- wire
			write                                               : in  std_logic                     := 'X';             -- wire
			frame_in                                            : out std_logic_vector(0 downto 0);                     -- wire
			eop                                                 : in  std_logic                     := 'X';             -- wire
			sop                                                 : in  std_logic                     := 'X';             -- wire
			Clock                                               : in  std_logic                     := 'X';             -- clk
			aclr                                                : in  std_logic                     := 'X';             -- reset
			valid                                               : in  std_logic                     := 'X';             -- wire
			row_counter                                         : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component Add_Frame_GN_Add_Frame_Add_Frame_Module;

	signal avalon_mm_slave_address_0_output_wire      : std_logic_vector(2 downto 0);  -- Avalon_MM_Slave_address_0:output -> Add_Frame_Add_Frame_Module_0:addr
	signal avalon_mm_slave_write_0_output_wire        : std_logic;                     -- Avalon_MM_Slave_write_0:output -> Add_Frame_Add_Frame_Module_0:write
	signal avalon_mm_slave_writedata_0_output_wire    : std_logic_vector(31 downto 0); -- Avalon_MM_Slave_writedata_0:output -> Add_Frame_Add_Frame_Module_0:writedata
	signal avalon_st_sink_data_0_output_wire          : std_logic_vector(23 downto 0); -- Avalon_ST_Sink_data_0:output -> Add_Frame_Add_Frame_Module_0:data_in
	signal avalon_st_sink_valid_0_output_wire         : std_logic;                     -- Avalon_ST_Sink_valid_0:output -> [Add_Frame_Add_Frame_Module_0:valid, Avalon_ST_Source_valid_0:input]
	signal avalon_st_sink_startofpacket_0_output_wire : std_logic;                     -- Avalon_ST_Sink_startofpacket_0:output -> [Add_Frame_Add_Frame_Module_0:sop, Avalon_ST_Source_startofpacket_0:input]
	signal avalon_st_sink_endofpacket_0_output_wire   : std_logic;                     -- Avalon_ST_Sink_endofpacket_0:output -> [Add_Frame_Add_Frame_Module_0:eop, Avalon_ST_Source_endofpacket_0:input]
	signal add_frame_add_frame_module_0_data_out_wire : std_logic_vector(23 downto 0); -- Add_Frame_Add_Frame_Module_0:data_out -> Avalon_ST_Source_data_0:input
	signal avalon_st_source_ready_0_output_wire       : std_logic;                     -- Avalon_ST_Source_ready_0:output -> Avalon_ST_Sink_ready_0:input
	signal clock_0_clock_output_reset                 : std_logic;                     -- Clock_0:aclr_out -> Add_Frame_Add_Frame_Module_0:aclr
	signal clock_0_clock_output_clk                   : std_logic;                     -- Clock_0:clock_out -> Add_Frame_Add_Frame_Module_0:Clock

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	avalon_mm_slave_address_0 : component alt_dspbuilder_port_GNS2GDLO5E
		port map (
			input  => Avalon_MM_Slave_address,               --  input.wire
			output => avalon_mm_slave_address_0_output_wire  -- output.wire
		);

	avalon_st_source_valid_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => avalon_st_sink_valid_0_output_wire, --  input.wire
			output => Avalon_ST_Source_valid              -- output.wire
		);

	avalon_mm_slave_writedata_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => Avalon_MM_Slave_writedata,               --  input.wire
			output => avalon_mm_slave_writedata_0_output_wire  -- output.wire
		);

	avalon_st_source_endofpacket_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => avalon_st_sink_endofpacket_0_output_wire, --  input.wire
			output => Avalon_ST_Source_endofpacket              -- output.wire
		);

	avalon_st_source_startofpacket_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => avalon_st_sink_startofpacket_0_output_wire, --  input.wire
			output => Avalon_ST_Source_startofpacket              -- output.wire
		);

	avalon_mm_slave_write_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Avalon_MM_Slave_write,               --  input.wire
			output => avalon_mm_slave_write_0_output_wire  -- output.wire
		);

	avalon_st_sink_data_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => Avalon_ST_Sink_data,               --  input.wire
			output => avalon_st_sink_data_0_output_wire  -- output.wire
		);

	avalon_st_sink_ready_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => avalon_st_source_ready_0_output_wire, --  input.wire
			output => Avalon_ST_Sink_ready                  -- output.wire
		);

	avalon_st_sink_startofpacket_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Avalon_ST_Sink_startofpacket,               --  input.wire
			output => avalon_st_sink_startofpacket_0_output_wire  -- output.wire
		);

	avalon_st_sink_endofpacket_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Avalon_ST_Sink_endofpacket,               --  input.wire
			output => avalon_st_sink_endofpacket_0_output_wire  -- output.wire
		);

	avalon_st_source_data_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => add_frame_add_frame_module_0_data_out_wire, --  input.wire
			output => Avalon_ST_Source_data                       -- output.wire
		);

	avalon_st_sink_valid_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Avalon_ST_Sink_valid,               --  input.wire
			output => avalon_st_sink_valid_0_output_wire  -- output.wire
		);

	add_frame_add_frame_module_0 : component Add_Frame_GN_Add_Frame_Add_Frame_Module
		port map (
			state                                               => Add_Frame_Add_Frame_Module_state,                    --                                               state.wire
			writedata                                           => avalon_mm_slave_writedata_0_output_wire,             --                                           writedata.wire
			Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_col => Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_col, -- Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_col.wire
			addr                                                => avalon_mm_slave_address_0_output_wire,               --                                                addr.wire
			data_in                                             => avalon_st_sink_data_0_output_wire,                   --                                             data_in.wire
			data_out                                            => add_frame_add_frame_module_0_data_out_wire,          --                                            data_out.wire
			Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_row => Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_row, -- Add_Frame_Add_Frame_Module_CTRL_DECODER_decoder_row.wire
			col_counter                                         => Add_Frame_Add_Frame_Module_col_counter,              --                                         col_counter.wire
			write                                               => avalon_mm_slave_write_0_output_wire,                 --                                               write.wire
			frame_in                                            => Add_Frame_Add_Frame_Module_frame_in,                 --                                            frame_in.wire
			eop                                                 => avalon_st_sink_endofpacket_0_output_wire,            --                                                 eop.wire
			sop                                                 => avalon_st_sink_startofpacket_0_output_wire,          --                                                 sop.wire
			Clock                                               => clock_0_clock_output_clk,                            --                                               Clock.clk
			aclr                                                => clock_0_clock_output_reset,                          --                                                    .reset
			valid                                               => avalon_st_sink_valid_0_output_wire,                  --                                               valid.wire
			row_counter                                         => Add_Frame_Add_Frame_Module_row_counter               --                                         row_counter.wire
		);

	avalon_st_source_ready_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Avalon_ST_Source_ready,               --  input.wire
			output => avalon_st_source_ready_0_output_wire  -- output.wire
		);

end architecture rtl; -- of Add_Frame_GN
