-- Add_Frame_GN_Add_Frame_Add_Frame_Module_Frame_Par.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.26.17:32:01

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Add_Frame_GN_Add_Frame_Add_Frame_Module_Frame_Par is
	port (
		vertex_col : out std_logic_vector(15 downto 0);                    -- vertex_col.wire
		vertex_row : out std_logic_vector(15 downto 0);                    -- vertex_row.wire
		Clock      : in  std_logic                     := '0';             --      Clock.clk
		aclr       : in  std_logic                     := '0';             --           .reset
		width      : out std_logic_vector(15 downto 0);                    --      width.wire
		data       : in  std_logic_vector(23 downto 0) := (others => '0'); --       data.wire
		writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --  writedata.wire
		write      : in  std_logic                     := '0';             --      write.wire
		height     : out std_logic_vector(15 downto 0);                    --     height.wire
		addr       : in  std_logic_vector(2 downto 0)  := (others => '0'); --       addr.wire
		sop        : in  std_logic                     := '0'              --        sop.wire
	);
end entity Add_Frame_GN_Add_Frame_Add_Frame_Module_Frame_Par;

architecture rtl of Add_Frame_GN_Add_Frame_Add_Frame_Module_Frame_Par is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_cast_GNNZHXLS76 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNNZHXLS76;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_port_GNS2GDLO5E is
		port (
			input  : in  std_logic_vector(2 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(2 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNS2GDLO5E;

	component alt_dspbuilder_port_GNBO6OMO5Y is
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNBO6OMO5Y;

	component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_decoder_GNBHXAVAPH is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNBHXAVAPH;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_decoder_GNSCEXJCJK is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNSCEXJCJK;

	component alt_dspbuilder_delay_GNKM23YKPN is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNKM23YKPN;

	component alt_dspbuilder_delay_GNC4JNSRBA is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNC4JNSRBA;

	component alt_dspbuilder_delay_GNH6PQLQQ2 is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNH6PQLQQ2;

	component alt_dspbuilder_decoder_GNQPHUITBS is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNQPHUITBS;

	component alt_dspbuilder_decoder_GN7W55JURN is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GN7W55JURN;

	component alt_dspbuilder_decoder_GNBT6YIKS3 is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNBT6YIKS3;

	signal decoder2sclrgnd_output_wire       : std_logic;                     -- Decoder2sclrGND:output -> Decoder2:sclr
	signal decoder2enavcc_output_wire        : std_logic;                     -- Decoder2enaVCC:output -> Decoder2:ena
	signal decoder3sclrgnd_output_wire       : std_logic;                     -- Decoder3sclrGND:output -> Decoder3:sclr
	signal decoder3enavcc_output_wire        : std_logic;                     -- Decoder3enaVCC:output -> Decoder3:ena
	signal decoder1sclrgnd_output_wire       : std_logic;                     -- Decoder1sclrGND:output -> Decoder1:sclr
	signal decoder1enavcc_output_wire        : std_logic;                     -- Decoder1enaVCC:output -> Decoder1:ena
	signal delay6sclrgnd_output_wire         : std_logic;                     -- Delay6sclrGND:output -> Delay6:sclr
	signal delay5sclrgnd_output_wire         : std_logic;                     -- Delay5sclrGND:output -> Delay5:sclr
	signal delay4sclrgnd_output_wire         : std_logic;                     -- Delay4sclrGND:output -> Delay4:sclr
	signal delay9sclrgnd_output_wire         : std_logic;                     -- Delay9sclrGND:output -> Delay9:sclr
	signal delay8sclrgnd_output_wire         : std_logic;                     -- Delay8sclrGND:output -> Delay8:sclr
	signal delay7sclrgnd_output_wire         : std_logic;                     -- Delay7sclrGND:output -> Delay7:sclr
	signal decoder7sclrgnd_output_wire       : std_logic;                     -- Decoder7sclrGND:output -> Decoder7:sclr
	signal decoder7enavcc_output_wire        : std_logic;                     -- Decoder7enaVCC:output -> Decoder7:ena
	signal delay10sclrgnd_output_wire        : std_logic;                     -- Delay10sclrGND:output -> Delay10:sclr
	signal decodersclrgnd_output_wire        : std_logic;                     -- DecodersclrGND:output -> Decoder:sclr
	signal decoderenavcc_output_wire         : std_logic;                     -- DecoderenaVCC:output -> Decoder:ena
	signal decoder6sclrgnd_output_wire       : std_logic;                     -- Decoder6sclrGND:output -> Decoder6:sclr
	signal decoder6enavcc_output_wire        : std_logic;                     -- Decoder6enaVCC:output -> Decoder6:ena
	signal delay11sclrgnd_output_wire        : std_logic;                     -- Delay11sclrGND:output -> Delay11:sclr
	signal decoder5sclrgnd_output_wire       : std_logic;                     -- Decoder5sclrGND:output -> Decoder5:sclr
	signal decoder5enavcc_output_wire        : std_logic;                     -- Decoder5enaVCC:output -> Decoder5:ena
	signal decoder4sclrgnd_output_wire       : std_logic;                     -- Decoder4sclrGND:output -> Decoder4:sclr
	signal decoder4enavcc_output_wire        : std_logic;                     -- Decoder4enaVCC:output -> Decoder4:ena
	signal writedata_0_output_wire           : std_logic_vector(31 downto 0); -- writedata_0:output -> [Bus_Conversion1:input, Bus_Conversion2:input, Bus_Conversion3:input, Bus_Conversion8:input]
	signal addr_0_output_wire                : std_logic_vector(2 downto 0);  -- addr_0:output -> [Decoder2:data, Decoder4:data, Decoder6:data, Decoder:data]
	signal bus_conversion8_output_wire       : std_logic_vector(15 downto 0); -- Bus_Conversion8:output -> Delay10:input
	signal delay10_output_wire               : std_logic_vector(15 downto 0); -- Delay10:output -> Delay11:input
	signal bus_conversion1_output_wire       : std_logic_vector(15 downto 0); -- Bus_Conversion1:output -> Delay4:input
	signal delay4_output_wire                : std_logic_vector(15 downto 0); -- Delay4:output -> Delay5:input
	signal bus_conversion2_output_wire       : std_logic_vector(15 downto 0); -- Bus_Conversion2:output -> Delay6:input
	signal delay6_output_wire                : std_logic_vector(15 downto 0); -- Delay6:output -> Delay7:input
	signal bus_conversion3_output_wire       : std_logic_vector(15 downto 0); -- Bus_Conversion3:output -> Delay8:input
	signal delay8_output_wire                : std_logic_vector(15 downto 0); -- Delay8:output -> Delay9:input
	signal data_0_output_wire                : std_logic_vector(23 downto 0); -- data_0:output -> [Decoder1:data, Decoder3:data, Decoder5:data, Decoder7:data]
	signal decoder_dec_wire                  : std_logic;                     -- Decoder:dec -> Logical_Bit_Operator1:data0
	signal write_0_output_wire               : std_logic;                     -- write_0:output -> [Logical_Bit_Operator1:data1, Logical_Bit_Operator4:data1, Logical_Bit_Operator6:data1, Logical_Bit_Operator8:data1]
	signal logical_bit_operator1_result_wire : std_logic;                     -- Logical_Bit_Operator1:result -> Delay4:ena
	signal sop_0_output_wire                 : std_logic;                     -- sop_0:output -> [Logical_Bit_Operator3:data0, Logical_Bit_Operator5:data0, Logical_Bit_Operator7:data0, Logical_Bit_Operator9:data0]
	signal decoder1_dec_wire                 : std_logic;                     -- Decoder1:dec -> Logical_Bit_Operator3:data1
	signal logical_bit_operator3_result_wire : std_logic;                     -- Logical_Bit_Operator3:result -> Delay5:ena
	signal decoder2_dec_wire                 : std_logic;                     -- Decoder2:dec -> Logical_Bit_Operator4:data0
	signal logical_bit_operator4_result_wire : std_logic;                     -- Logical_Bit_Operator4:result -> Delay6:ena
	signal decoder3_dec_wire                 : std_logic;                     -- Decoder3:dec -> Logical_Bit_Operator5:data1
	signal logical_bit_operator5_result_wire : std_logic;                     -- Logical_Bit_Operator5:result -> Delay7:ena
	signal decoder4_dec_wire                 : std_logic;                     -- Decoder4:dec -> Logical_Bit_Operator6:data0
	signal logical_bit_operator6_result_wire : std_logic;                     -- Logical_Bit_Operator6:result -> Delay8:ena
	signal decoder5_dec_wire                 : std_logic;                     -- Decoder5:dec -> Logical_Bit_Operator7:data1
	signal logical_bit_operator7_result_wire : std_logic;                     -- Logical_Bit_Operator7:result -> Delay9:ena
	signal decoder6_dec_wire                 : std_logic;                     -- Decoder6:dec -> Logical_Bit_Operator8:data0
	signal logical_bit_operator8_result_wire : std_logic;                     -- Logical_Bit_Operator8:result -> Delay10:ena
	signal decoder7_dec_wire                 : std_logic;                     -- Decoder7:dec -> Logical_Bit_Operator9:data1
	signal logical_bit_operator9_result_wire : std_logic;                     -- Logical_Bit_Operator9:result -> Delay11:ena
	signal delay5_output_wire                : std_logic_vector(15 downto 0); -- Delay5:output -> vertex_col_0:input
	signal delay7_output_wire                : std_logic_vector(15 downto 0); -- Delay7:output -> vertex_row_0:input
	signal delay9_output_wire                : std_logic_vector(15 downto 0); -- Delay9:output -> width_0:input
	signal delay11_output_wire               : std_logic_vector(15 downto 0); -- Delay11:output -> height_0:input
	signal clock_0_clock_output_reset        : std_logic;                     -- Clock_0:aclr_out -> [Decoder1:aclr, Decoder2:aclr, Decoder3:aclr, Decoder4:aclr, Decoder5:aclr, Decoder6:aclr, Decoder7:aclr, Decoder:aclr, Delay10:aclr, Delay11:aclr, Delay4:aclr, Delay5:aclr, Delay6:aclr, Delay7:aclr, Delay8:aclr, Delay9:aclr]
	signal clock_0_clock_output_clk          : std_logic;                     -- Clock_0:clock_out -> [Decoder1:clock, Decoder2:clock, Decoder3:clock, Decoder4:clock, Decoder5:clock, Decoder6:clock, Decoder7:clock, Decoder:clock, Delay10:clock, Delay11:clock, Delay4:clock, Delay5:clock, Delay6:clock, Delay7:clock, Delay8:clock, Delay9:clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	bus_conversion1 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => writedata_0_output_wire,     --  input.wire
			output => bus_conversion1_output_wire  -- output.wire
		);

	bus_conversion2 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => writedata_0_output_wire,     --  input.wire
			output => bus_conversion2_output_wire  -- output.wire
		);

	bus_conversion3 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => writedata_0_output_wire,     --  input.wire
			output => bus_conversion3_output_wire  -- output.wire
		);

	writedata_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => writedata,               --  input.wire
			output => writedata_0_output_wire  -- output.wire
		);

	data_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => data,               --  input.wire
			output => data_0_output_wire  -- output.wire
		);

	addr_0 : component alt_dspbuilder_port_GNS2GDLO5E
		port map (
			input  => addr,               --  input.wire
			output => addr_0_output_wire  -- output.wire
		);

	vertex_row_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => delay7_output_wire, --  input.wire
			output => vertex_row          -- output.wire
		);

	logical_bit_operator7 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator7_result_wire, -- result.wire
			data0  => sop_0_output_wire,                 --  data0.wire
			data1  => decoder5_dec_wire                  --  data1.wire
		);

	logical_bit_operator6 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator6_result_wire, -- result.wire
			data0  => decoder4_dec_wire,                 --  data0.wire
			data1  => write_0_output_wire                --  data1.wire
		);

	vertex_col_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => delay5_output_wire, --  input.wire
			output => vertex_col          -- output.wire
		);

	logical_bit_operator5 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator5_result_wire, -- result.wire
			data0  => sop_0_output_wire,                 --  data0.wire
			data1  => decoder3_dec_wire                  --  data1.wire
		);

	height_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => delay11_output_wire, --  input.wire
			output => height               -- output.wire
		);

	logical_bit_operator4 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator4_result_wire, -- result.wire
			data0  => decoder2_dec_wire,                 --  data0.wire
			data1  => write_0_output_wire                --  data1.wire
		);

	logical_bit_operator9 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator9_result_wire, -- result.wire
			data0  => sop_0_output_wire,                 --  data0.wire
			data1  => decoder7_dec_wire                  --  data1.wire
		);

	logical_bit_operator8 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator8_result_wire, -- result.wire
			data0  => decoder6_dec_wire,                 --  data0.wire
			data1  => write_0_output_wire                --  data1.wire
		);

	write_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => write,               --  input.wire
			output => write_0_output_wire  -- output.wire
		);

	logical_bit_operator3 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator3_result_wire, -- result.wire
			data0  => sop_0_output_wire,                 --  data0.wire
			data1  => decoder1_dec_wire                  --  data1.wire
		);

	logical_bit_operator1 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator1_result_wire, -- result.wire
			data0  => decoder_dec_wire,                  --  data0.wire
			data1  => write_0_output_wire                --  data1.wire
		);

	decoder2 : component alt_dspbuilder_decoder_GNBHXAVAPH
		generic map (
			decode   => "010",
			pipeline => 1,
			width    => 3
		)
		port map (
			clock => clock_0_clock_output_clk,    -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,  --           .reset
			data  => addr_0_output_wire,          --       data.wire
			dec   => decoder2_dec_wire,           --        dec.wire
			sclr  => decoder2sclrgnd_output_wire, --       sclr.wire
			ena   => decoder2enavcc_output_wire   --        ena.wire
		);

	decoder2sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder2sclrgnd_output_wire  -- output.wire
		);

	decoder2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder2enavcc_output_wire  -- output.wire
		);

	decoder3 : component alt_dspbuilder_decoder_GNSCEXJCJK
		generic map (
			decode   => "000000000000000000001111",
			pipeline => 0,
			width    => 24
		)
		port map (
			clock => clock_0_clock_output_clk,    -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,  --           .reset
			data  => data_0_output_wire,          --       data.wire
			dec   => decoder3_dec_wire,           --        dec.wire
			sclr  => decoder3sclrgnd_output_wire, --       sclr.wire
			ena   => decoder3enavcc_output_wire   --        ena.wire
		);

	decoder3sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder3sclrgnd_output_wire  -- output.wire
		);

	decoder3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder3enavcc_output_wire  -- output.wire
		);

	decoder1 : component alt_dspbuilder_decoder_GNSCEXJCJK
		generic map (
			decode   => "000000000000000000001111",
			pipeline => 0,
			width    => 24
		)
		port map (
			clock => clock_0_clock_output_clk,    -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,  --           .reset
			data  => data_0_output_wire,          --       data.wire
			dec   => decoder1_dec_wire,           --        dec.wire
			sclr  => decoder1sclrgnd_output_wire, --       sclr.wire
			ena   => decoder1enavcc_output_wire   --        ena.wire
		);

	decoder1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder1sclrgnd_output_wire  -- output.wire
		);

	decoder1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder1enavcc_output_wire  -- output.wire
		);

	width_0 : component alt_dspbuilder_port_GNBO6OMO5Y
		port map (
			input  => delay9_output_wire, --  input.wire
			output => width               -- output.wire
		);

	delay6 : component alt_dspbuilder_delay_GNKM23YKPN
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0000000001100100",
			width      => 16
		)
		port map (
			input  => bus_conversion2_output_wire,       --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay6_output_wire,                --     output.wire
			sclr   => delay6sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator4_result_wire  --        ena.wire
		);

	delay6sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay6sclrgnd_output_wire  -- output.wire
		);

	delay5 : component alt_dspbuilder_delay_GNC4JNSRBA
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0000000100101100",
			width      => 16
		)
		port map (
			input  => delay4_output_wire,                --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay5_output_wire,                --     output.wire
			sclr   => delay5sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator3_result_wire  --        ena.wire
		);

	delay5sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay5sclrgnd_output_wire  -- output.wire
		);

	delay4 : component alt_dspbuilder_delay_GNC4JNSRBA
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0000000100101100",
			width      => 16
		)
		port map (
			input  => bus_conversion1_output_wire,       --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay4_output_wire,                --     output.wire
			sclr   => delay4sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator1_result_wire  --        ena.wire
		);

	delay4sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay4sclrgnd_output_wire  -- output.wire
		);

	sop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sop,               --  input.wire
			output => sop_0_output_wire  -- output.wire
		);

	delay9 : component alt_dspbuilder_delay_GNH6PQLQQ2
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0000000000110010",
			width      => 16
		)
		port map (
			input  => delay8_output_wire,                --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay9_output_wire,                --     output.wire
			sclr   => delay9sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator7_result_wire  --        ena.wire
		);

	delay9sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay9sclrgnd_output_wire  -- output.wire
		);

	delay8 : component alt_dspbuilder_delay_GNH6PQLQQ2
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0000000000110010",
			width      => 16
		)
		port map (
			input  => bus_conversion3_output_wire,       --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay8_output_wire,                --     output.wire
			sclr   => delay8sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator6_result_wire  --        ena.wire
		);

	delay8sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay8sclrgnd_output_wire  -- output.wire
		);

	delay7 : component alt_dspbuilder_delay_GNKM23YKPN
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0000000001100100",
			width      => 16
		)
		port map (
			input  => delay6_output_wire,                --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay7_output_wire,                --     output.wire
			sclr   => delay7sclrgnd_output_wire,         --       sclr.wire
			ena    => logical_bit_operator5_result_wire  --        ena.wire
		);

	delay7sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay7sclrgnd_output_wire  -- output.wire
		);

	bus_conversion8 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => writedata_0_output_wire,     --  input.wire
			output => bus_conversion8_output_wire  -- output.wire
		);

	decoder7 : component alt_dspbuilder_decoder_GNSCEXJCJK
		generic map (
			decode   => "000000000000000000001111",
			pipeline => 0,
			width    => 24
		)
		port map (
			clock => clock_0_clock_output_clk,    -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,  --           .reset
			data  => data_0_output_wire,          --       data.wire
			dec   => decoder7_dec_wire,           --        dec.wire
			sclr  => decoder7sclrgnd_output_wire, --       sclr.wire
			ena   => decoder7enavcc_output_wire   --        ena.wire
		);

	decoder7sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder7sclrgnd_output_wire  -- output.wire
		);

	decoder7enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder7enavcc_output_wire  -- output.wire
		);

	delay10 : component alt_dspbuilder_delay_GNC4JNSRBA
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0000000100101100",
			width      => 16
		)
		port map (
			input  => bus_conversion8_output_wire,       --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay10_output_wire,               --     output.wire
			sclr   => delay10sclrgnd_output_wire,        --       sclr.wire
			ena    => logical_bit_operator8_result_wire  --        ena.wire
		);

	delay10sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay10sclrgnd_output_wire  -- output.wire
		);

	decoder : component alt_dspbuilder_decoder_GNQPHUITBS
		generic map (
			decode   => "001",
			pipeline => 1,
			width    => 3
		)
		port map (
			clock => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset, --           .reset
			data  => addr_0_output_wire,         --       data.wire
			dec   => decoder_dec_wire,           --        dec.wire
			sclr  => decodersclrgnd_output_wire, --       sclr.wire
			ena   => decoderenavcc_output_wire   --        ena.wire
		);

	decodersclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decodersclrgnd_output_wire  -- output.wire
		);

	decoderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoderenavcc_output_wire  -- output.wire
		);

	decoder6 : component alt_dspbuilder_decoder_GN7W55JURN
		generic map (
			decode   => "100",
			pipeline => 1,
			width    => 3
		)
		port map (
			clock => clock_0_clock_output_clk,    -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,  --           .reset
			data  => addr_0_output_wire,          --       data.wire
			dec   => decoder6_dec_wire,           --        dec.wire
			sclr  => decoder6sclrgnd_output_wire, --       sclr.wire
			ena   => decoder6enavcc_output_wire   --        ena.wire
		);

	decoder6sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder6sclrgnd_output_wire  -- output.wire
		);

	decoder6enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder6enavcc_output_wire  -- output.wire
		);

	delay11 : component alt_dspbuilder_delay_GNC4JNSRBA
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0000000100101100",
			width      => 16
		)
		port map (
			input  => delay10_output_wire,               --      input.wire
			clock  => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,        --           .reset
			output => delay11_output_wire,               --     output.wire
			sclr   => delay11sclrgnd_output_wire,        --       sclr.wire
			ena    => logical_bit_operator9_result_wire  --        ena.wire
		);

	delay11sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay11sclrgnd_output_wire  -- output.wire
		);

	decoder5 : component alt_dspbuilder_decoder_GNSCEXJCJK
		generic map (
			decode   => "000000000000000000001111",
			pipeline => 0,
			width    => 24
		)
		port map (
			clock => clock_0_clock_output_clk,    -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,  --           .reset
			data  => data_0_output_wire,          --       data.wire
			dec   => decoder5_dec_wire,           --        dec.wire
			sclr  => decoder5sclrgnd_output_wire, --       sclr.wire
			ena   => decoder5enavcc_output_wire   --        ena.wire
		);

	decoder5sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder5sclrgnd_output_wire  -- output.wire
		);

	decoder5enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder5enavcc_output_wire  -- output.wire
		);

	decoder4 : component alt_dspbuilder_decoder_GNBT6YIKS3
		generic map (
			decode   => "011",
			pipeline => 1,
			width    => 3
		)
		port map (
			clock => clock_0_clock_output_clk,    -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,  --           .reset
			data  => addr_0_output_wire,          --       data.wire
			dec   => decoder4_dec_wire,           --        dec.wire
			sclr  => decoder4sclrgnd_output_wire, --       sclr.wire
			ena   => decoder4enavcc_output_wire   --        ena.wire
		);

	decoder4sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder4sclrgnd_output_wire  -- output.wire
		);

	decoder4enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder4enavcc_output_wire  -- output.wire
		);

end architecture rtl; -- of Add_Frame_GN_Add_Frame_Add_Frame_Module_Frame_Par
