-- Add_Frame_GN_Add_Frame_Add_Frame_Module.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.27.11:15:10

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Add_Frame_GN_Add_Frame_Add_Frame_Module is
	port (
		data_out  : out std_logic_vector(23 downto 0);                    --  data_out.wire
		addr      : in  std_logic_vector(2 downto 0)  := (others => '0'); --      addr.wire
		write     : in  std_logic                     := '0';             --     write.wire
		writedata : in  std_logic_vector(31 downto 0) := (others => '0'); -- writedata.wire
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		aclr      : in  std_logic                     := '0';             --          .reset
		sop       : in  std_logic                     := '0';             --       sop.wire
		eop       : in  std_logic                     := '0';             --       eop.wire
		valid     : in  std_logic                     := '0';             --     valid.wire
		data_in   : in  std_logic_vector(23 downto 0) := (others => '0')  --   data_in.wire
	);
end entity Add_Frame_GN_Add_Frame_Add_Frame_Module;

architecture rtl of Add_Frame_GN_Add_Frame_Add_Frame_Module is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_pipelined_adder_GNWEIMU3MK is
		generic (
			width    : natural := 0;
			pipeline : integer := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNWEIMU3MK;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_pipelined_adder_GNTWZRTG4I is
		generic (
			width    : natural := 0;
			pipeline : integer := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNTWZRTG4I;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_constant_GNWFCSDEFM is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(15 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNWFCSDEFM;

	component alt_dspbuilder_constant_GNLMV7GZFA is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNLMV7GZFA;

	component alt_dspbuilder_port_GNS2GDLO5E is
		port (
			input  : in  std_logic_vector(2 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(2 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNS2GDLO5E;

	component alt_dspbuilder_constant_GNZEH3JAKA is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNZEH3JAKA;

	component alt_dspbuilder_constant_GNNKZSYI73 is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNNKZSYI73;

	component alt_dspbuilder_constant_GNGITJD4MB is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNGITJD4MB;

	component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V;

	component alt_dspbuilder_logical_bit_op_GN5A3KLAEC is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'; -- wire
			data2  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GN5A3KLAEC;

	component alt_dspbuilder_logical_bit_op_GNKUBZL4TE is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNKUBZL4TE;

	component alt_dspbuilder_logical_bit_op_GNUQ2R64DV is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNUQ2R64DV;

	component alt_dspbuilder_constant_GNNTMI25OE is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNNTMI25OE;

	component alt_dspbuilder_constant_GNIJTURCWG is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNIJTURCWG;

	component alt_dspbuilder_if_statement_GNHRNNRV37 is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			c    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			d    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			e    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			f    : in  std_logic_vector(15 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNHRNNRV37;

	component Add_Frame_GN_Add_Frame_Add_Frame_Module_FRAME_PARAMETER is
		port (
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			data       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			height     : out std_logic_vector(15 downto 0);                    -- wire
			Clock      : in  std_logic                     := 'X';             -- clk
			aclr       : in  std_logic                     := 'X';             -- reset
			write      : in  std_logic                     := 'X';             -- wire
			width      : out std_logic_vector(15 downto 0);                    -- wire
			sop        : in  std_logic                     := 'X';             -- wire
			enble      : out std_logic_vector(0 downto 0);                     -- wire
			addr       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- wire
			color      : out std_logic_vector(2 downto 0);                     -- wire
			vertex_col : out std_logic_vector(15 downto 0);                    -- wire
			vertex_row : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component Add_Frame_GN_Add_Frame_Add_Frame_Module_FRAME_PARAMETER;

	component Add_Frame_GN_Add_Frame_Add_Frame_Module_CTRL_DECODER is
		port (
			height : out std_logic_vector(15 downto 0);                    -- wire
			width  : out std_logic_vector(15 downto 0);                    -- wire
			sop    : in  std_logic                     := 'X';             -- wire
			Clock  : in  std_logic                     := 'X';             -- clk
			aclr   : in  std_logic                     := 'X';             -- reset
			data   : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			valid  : in  std_logic                     := 'X'              -- wire
		);
	end component Add_Frame_GN_Add_Frame_Add_Frame_Module_CTRL_DECODER;

	component alt_dspbuilder_single_pulse_GN2XGKTRR3 is
		generic (
			delay         : positive := 1;
			signal_type   : string   := "Impulse";
			impulse_width : positive := 1
		);
		port (
			aclr   : in  std_logic := 'X'; -- clk
			clock  : in  std_logic := 'X'; -- clk
			ena    : in  std_logic := 'X'; -- wire
			result : out std_logic;        -- wire
			sclr   : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_single_pulse_GN2XGKTRR3;

	component alt_dspbuilder_if_statement_GNUCFELPE2 is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(15 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNUCFELPE2;

	component alt_dspbuilder_counter_GNCXSYJEM5 is
		generic (
			use_usr_aclr : string  := "false";
			use_ena      : string  := "false";
			use_cin      : string  := "false";
			use_sset     : string  := "false";
			ndirection   : natural := 1;
			svalue       : string  := "0";
			use_sload    : string  := "false";
			use_sclr     : string  := "false";
			use_cout     : string  := "false";
			modulus      : integer := 256;
			use_cnt_ena  : string  := "false";
			width        : natural := 8;
			use_aset     : string  := "false";
			use_aload    : string  := "false";
			avalue       : string  := "0"
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			aload     : in  std_logic                          := 'X';             -- wire
			aset      : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cnt_ena   : in  std_logic                          := 'X';             -- wire
			cout      : out std_logic;                                             -- wire
			data      : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			direction : in  std_logic                          := 'X';             -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			q         : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr      : in  std_logic                          := 'X';             -- wire
			sload     : in  std_logic                          := 'X';             -- wire
			sset      : in  std_logic                          := 'X';             -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_counter_GNCXSYJEM5;

	component alt_dspbuilder_if_statement_GN7VA7SRUP is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			c    : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GN7VA7SRUP;

	component FrameControl is
		port (
			clock    : in  std_logic                    := 'X'; -- clk
			ctrl_in  : in  std_logic                    := 'X'; -- wire
			data_in  : in  std_logic                    := 'X'; -- wire
			frame_in : in  std_logic                    := 'X'; -- wire
			reset    : in  std_logic                    := 'X'; -- wire
			state    : out std_logic_vector(2 downto 0)         -- wire
		);
	end component FrameControl;

	component alt_dspbuilder_delay_GNHYCSAEGT is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNHYCSAEGT;

	component alt_dspbuilder_multiplexer_GNRF25WCVA is
		generic (
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0;
			width                  : positive := 8;
			pipeline               : natural  := 0;
			number_inputs          : natural  := 4
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(23 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in2       : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNRF25WCVA;

	component alt_dspbuilder_delay_GNUECIBFDH is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNUECIBFDH;

	component alt_dspbuilder_multiplexer_GNHHROOGAI is
		generic (
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0;
			width                  : positive := 8;
			pipeline               : natural  := 0;
			number_inputs          : natural  := 4
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(23 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in2       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in3       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in4       : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNHHROOGAI;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_cast_GNSB3OXIQS is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			output : out std_logic                                        -- wire
		);
	end component alt_dspbuilder_cast_GNSB3OXIQS;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	component alt_dspbuilder_cast_GNLWRZWTQF is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(2 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(2 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNLWRZWTQF;

	signal pipelined_adder3user_aclrgnd_output_wire                     : std_logic;                     -- Pipelined_Adder3user_aclrGND:output -> Pipelined_Adder3:user_aclr
	signal pipelined_adder3enavcc_output_wire                           : std_logic;                     -- Pipelined_Adder3enaVCC:output -> Pipelined_Adder3:ena
	signal pipelined_adder4user_aclrgnd_output_wire                     : std_logic;                     -- Pipelined_Adder4user_aclrGND:output -> Pipelined_Adder4:user_aclr
	signal pipelined_adder4enavcc_output_wire                           : std_logic;                     -- Pipelined_Adder4enaVCC:output -> Pipelined_Adder4:ena
	signal pipelined_adder1user_aclrgnd_output_wire                     : std_logic;                     -- Pipelined_Adder1user_aclrGND:output -> Pipelined_Adder1:user_aclr
	signal pipelined_adder1enavcc_output_wire                           : std_logic;                     -- Pipelined_Adder1enaVCC:output -> Pipelined_Adder1:ena
	signal pipelined_adder2user_aclrgnd_output_wire                     : std_logic;                     -- Pipelined_Adder2user_aclrGND:output -> Pipelined_Adder2:user_aclr
	signal pipelined_adder2enavcc_output_wire                           : std_logic;                     -- Pipelined_Adder2enaVCC:output -> Pipelined_Adder2:ena
	signal single_pulsesclrgnd_output_wire                              : std_logic;                     -- Single_PulsesclrGND:output -> Single_Pulse:sclr
	signal single_pulseenavcc_output_wire                               : std_logic;                     -- Single_PulseenaVCC:output -> Single_Pulse:ena
	signal pipelined_adderuser_aclrgnd_output_wire                      : std_logic;                     -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal pipelined_adderenavcc_output_wire                            : std_logic;                     -- Pipelined_AdderenaVCC:output -> Pipelined_Adder:ena
	signal delay3sclrgnd_output_wire                                    : std_logic;                     -- Delay3sclrGND:output -> Delay3:sclr
	signal delay3enavcc_output_wire                                     : std_logic;                     -- Delay3enaVCC:output -> Delay3:ena
	signal multiplexer1user_aclrgnd_output_wire                         : std_logic;                     -- Multiplexer1user_aclrGND:output -> Multiplexer1:user_aclr
	signal multiplexer1enavcc_output_wire                               : std_logic;                     -- Multiplexer1enaVCC:output -> Multiplexer1:ena
	signal multiplexer2user_aclrgnd_output_wire                         : std_logic;                     -- Multiplexer2user_aclrGND:output -> Multiplexer2:user_aclr
	signal multiplexer2enavcc_output_wire                               : std_logic;                     -- Multiplexer2enaVCC:output -> Multiplexer2:ena
	signal delay2sclrgnd_output_wire                                    : std_logic;                     -- Delay2sclrGND:output -> Delay2:sclr
	signal delay2enavcc_output_wire                                     : std_logic;                     -- Delay2enaVCC:output -> Delay2:ena
	signal sop_0_output_wire                                            : std_logic;                     -- sop_0:output -> [Add_Frame_Add_Frame_Module_CTRL_DECODER_0:sop, Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:sop, Logical_Bit_Operator:data1]
	signal valid_0_output_wire                                          : std_logic;                     -- valid_0:output -> [Add_Frame_Add_Frame_Module_CTRL_DECODER_0:valid, Logical_Bit_Operator1:data1, Logical_Bit_Operator6:data2]
	signal delay3_output_wire                                           : std_logic_vector(0 downto 0);  -- Delay3:output -> [Delay1:input, cast10:input]
	signal addr_0_output_wire                                           : std_logic_vector(2 downto 0);  -- addr_0:output -> Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:addr
	signal write_0_output_wire                                          : std_logic;                     -- write_0:output -> Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:write
	signal writedata_0_output_wire                                      : std_logic_vector(31 downto 0); -- writedata_0:output -> Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:writedata
	signal data_in_0_output_wire                                        : std_logic_vector(23 downto 0); -- data_in_0:output -> [Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:data, If_Statement1:a, Multiplexer1:in0, Multiplexer1:in1]
	signal counter_q_wire                                               : std_logic_vector(15 downto 0); -- Counter:q -> [If_Statement2:b, If_Statement3:b, If_Statement:a]
	signal add_frame_add_frame_module_frame_parameter_0_vertex_col_wire : std_logic_vector(15 downto 0); -- Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:vertex_col -> [If_Statement:b, Pipelined_Adder:dataa]
	signal counter1_q_wire                                              : std_logic_vector(15 downto 0); -- Counter1:q -> [If_Statement4:b, If_Statement:d]
	signal add_frame_add_frame_module_frame_parameter_0_vertex_row_wire : std_logic_vector(15 downto 0); -- Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:vertex_row -> [If_Statement:e, Pipelined_Adder1:dataa]
	signal constant3_output_wire                                        : std_logic_vector(23 downto 0); -- Constant3:output -> If_Statement1:b
	signal constant4_output_wire                                        : std_logic_vector(23 downto 0); -- Constant4:output -> If_Statement1:c
	signal if_statement1_true_wire                                      : std_logic;                     -- If_Statement1:true -> Logical_Bit_Operator:data0
	signal logical_bit_operator1_result_wire                            : std_logic;                     -- Logical_Bit_Operator1:result -> Counter:cnt_ena
	signal eop_0_output_wire                                            : std_logic;                     -- eop_0:output -> Logical_Bit_Operator2:data0
	signal logical_bit_operator3_result_wire                            : std_logic;                     -- Logical_Bit_Operator3:result -> Frame_Control:ctrl_in
	signal if_statement4_true_wire                                      : std_logic;                     -- If_Statement4:true -> Logical_Bit_Operator4:data0
	signal if_statement3_true_wire                                      : std_logic;                     -- If_Statement3:true -> Logical_Bit_Operator4:data1
	signal logical_bit_operator4_result_wire                            : std_logic;                     -- Logical_Bit_Operator4:result -> Counter:sclr
	signal logical_bit_operator5_result_wire                            : std_logic;                     -- Logical_Bit_Operator5:result -> Counter1:sclr
	signal if_statement2_true_wire                                      : std_logic;                     -- If_Statement2:true -> Logical_Bit_Operator6:data1
	signal logical_bit_operator6_result_wire                            : std_logic;                     -- Logical_Bit_Operator6:result -> Counter1:cnt_ena
	signal if_statement_true_wire                                       : std_logic;                     -- If_Statement:true -> Logical_Bit_Operator7:data1
	signal logical_bit_operator7_result_wire                            : std_logic;                     -- Logical_Bit_Operator7:result -> Frame_Control:frame_in
	signal multiplexer1_result_wire                                     : std_logic_vector(23 downto 0); -- Multiplexer1:result -> [Add_Frame_Add_Frame_Module_CTRL_DECODER_0:data, data_out_0:input]
	signal add_frame_add_frame_module_frame_parameter_0_color_wire      : std_logic_vector(2 downto 0);  -- Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:color -> Multiplexer2:sel
	signal constant5_output_wire                                        : std_logic_vector(23 downto 0); -- Constant5:output -> Multiplexer2:in0
	signal constant7_output_wire                                        : std_logic_vector(23 downto 0); -- Constant7:output -> Multiplexer2:in1
	signal constant9_output_wire                                        : std_logic_vector(23 downto 0); -- Constant9:output -> Multiplexer2:in2
	signal constant10_output_wire                                       : std_logic_vector(23 downto 0); -- Constant10:output -> Multiplexer2:in3
	signal constant11_output_wire                                       : std_logic_vector(23 downto 0); -- Constant11:output -> Multiplexer2:in4
	signal multiplexer2_result_wire                                     : std_logic_vector(23 downto 0); -- Multiplexer2:result -> Multiplexer1:in2
	signal add_frame_add_frame_module_frame_parameter_0_width_wire      : std_logic_vector(15 downto 0); -- Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:width -> Pipelined_Adder:datab
	signal pipelined_adder_result_wire                                  : std_logic_vector(15 downto 0); -- Pipelined_Adder:result -> If_Statement:c
	signal add_frame_add_frame_module_frame_parameter_0_height_wire     : std_logic_vector(15 downto 0); -- Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:height -> Pipelined_Adder1:datab
	signal pipelined_adder1_result_wire                                 : std_logic_vector(15 downto 0); -- Pipelined_Adder1:result -> If_Statement:f
	signal constant1_output_wire                                        : std_logic_vector(15 downto 0); -- Constant1:output -> Pipelined_Adder2:datab
	signal pipelined_adder2_result_wire                                 : std_logic_vector(15 downto 0); -- Pipelined_Adder2:result -> If_Statement2:a
	signal add_frame_add_frame_module_ctrl_decoder_0_width_wire         : std_logic_vector(15 downto 0); -- Add_Frame_Add_Frame_Module_CTRL_DECODER_0:width -> Pipelined_Adder3:dataa
	signal constant6_output_wire                                        : std_logic_vector(15 downto 0); -- Constant6:output -> Pipelined_Adder3:datab
	signal pipelined_adder3_result_wire                                 : std_logic_vector(15 downto 0); -- Pipelined_Adder3:result -> [If_Statement3:a, Pipelined_Adder2:dataa]
	signal add_frame_add_frame_module_ctrl_decoder_0_height_wire        : std_logic_vector(15 downto 0); -- Add_Frame_Add_Frame_Module_CTRL_DECODER_0:height -> Pipelined_Adder4:dataa
	signal constant8_output_wire                                        : std_logic_vector(15 downto 0); -- Constant8:output -> Pipelined_Adder4:datab
	signal pipelined_adder4_result_wire                                 : std_logic_vector(15 downto 0); -- Pipelined_Adder4:result -> If_Statement4:a
	signal single_pulse_result_wire                                     : std_logic;                     -- Single_Pulse:result -> Frame_Control:reset
	signal delay2_output_wire                                           : std_logic_vector(0 downto 0);  -- Delay2:output -> cast9:input
	signal cast9_output_wire                                            : std_logic;                     -- cast9:output -> Delay1:sclr
	signal cast10_output_wire                                           : std_logic;                     -- cast10:output -> Delay1:ena
	signal delay1_output_wire                                           : std_logic_vector(0 downto 0);  -- Delay1:output -> [cast11:input, cast13:input, cast14:input, cast16:input, cast17:input, cast18:input]
	signal cast11_output_wire                                           : std_logic;                     -- cast11:output -> Frame_Control:data_in
	signal logical_bit_operator_result_wire                             : std_logic;                     -- Logical_Bit_Operator:result -> cast12:input
	signal cast12_output_wire                                           : std_logic_vector(0 downto 0);  -- cast12:output -> Delay3:input
	signal cast13_output_wire                                           : std_logic;                     -- cast13:output -> Logical_Bit_Operator1:data0
	signal cast14_output_wire                                           : std_logic;                     -- cast14:output -> Logical_Bit_Operator2:data1
	signal logical_bit_operator2_result_wire                            : std_logic;                     -- Logical_Bit_Operator2:result -> cast15:input
	signal cast15_output_wire                                           : std_logic_vector(0 downto 0);  -- cast15:output -> Delay2:input
	signal cast16_output_wire                                           : std_logic;                     -- cast16:output -> Logical_Bit_Operator3:data0
	signal cast17_output_wire                                           : std_logic;                     -- cast17:output -> Logical_Bit_Operator5:data0
	signal cast18_output_wire                                           : std_logic;                     -- cast18:output -> Logical_Bit_Operator6:data0
	signal add_frame_add_frame_module_frame_parameter_0_enble_wire      : std_logic_vector(0 downto 0);  -- Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:enble -> cast19:input
	signal cast19_output_wire                                           : std_logic;                     -- cast19:output -> Logical_Bit_Operator7:data0
	signal frame_control_state_wire                                     : std_logic_vector(2 downto 0);  -- Frame_Control:state -> cast20:input
	signal cast20_output_wire                                           : std_logic_vector(2 downto 0);  -- cast20:output -> Multiplexer1:sel
	signal clock_0_clock_output_reset                                   : std_logic;                     -- Clock_0:aclr_out -> [Add_Frame_Add_Frame_Module_CTRL_DECODER_0:aclr, Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:aclr, Counter1:aclr, Counter:aclr, Delay1:aclr, Delay2:aclr, Delay3:aclr, Multiplexer1:aclr, Multiplexer2:aclr, Pipelined_Adder1:aclr, Pipelined_Adder2:aclr, Pipelined_Adder3:aclr, Pipelined_Adder4:aclr, Pipelined_Adder:aclr, Single_Pulse:aclr]
	signal clock_0_clock_output_clk                                     : std_logic;                     -- Clock_0:clock_out -> [Add_Frame_Add_Frame_Module_CTRL_DECODER_0:Clock, Add_Frame_Add_Frame_Module_FRAME_PARAMETER_0:Clock, Counter1:clock, Counter:clock, Delay1:clock, Delay2:clock, Delay3:clock, Frame_Control:clock, Multiplexer1:clock, Multiplexer2:clock, Pipelined_Adder1:clock, Pipelined_Adder2:clock, Pipelined_Adder3:clock, Pipelined_Adder4:clock, Pipelined_Adder:clock, Single_Pulse:clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	pipelined_adder3 : component alt_dspbuilder_pipelined_adder_GNWEIMU3MK
		generic map (
			width    => 16,
			pipeline => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,                             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                           --           .reset
			dataa     => add_frame_add_frame_module_ctrl_decoder_0_width_wire, --      dataa.wire
			datab     => constant6_output_wire,                                --      datab.wire
			result    => pipelined_adder3_result_wire,                         --     result.wire
			user_aclr => pipelined_adder3user_aclrgnd_output_wire,             --  user_aclr.wire
			ena       => pipelined_adder3enavcc_output_wire                    --        ena.wire
		);

	pipelined_adder3user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder3user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder3enavcc_output_wire  -- output.wire
		);

	pipelined_adder4 : component alt_dspbuilder_pipelined_adder_GNWEIMU3MK
		generic map (
			width    => 16,
			pipeline => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,                              -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                            --           .reset
			dataa     => add_frame_add_frame_module_ctrl_decoder_0_height_wire, --      dataa.wire
			datab     => constant8_output_wire,                                 --      datab.wire
			result    => pipelined_adder4_result_wire,                          --     result.wire
			user_aclr => pipelined_adder4user_aclrgnd_output_wire,              --  user_aclr.wire
			ena       => pipelined_adder4enavcc_output_wire                     --        ena.wire
		);

	pipelined_adder4user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder4user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder4enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder4enavcc_output_wire  -- output.wire
		);

	valid_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => valid,               --  input.wire
			output => valid_0_output_wire  -- output.wire
		);

	pipelined_adder1 : component alt_dspbuilder_pipelined_adder_GNTWZRTG4I
		generic map (
			width    => 16,
			pipeline => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,                                     -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                                   --           .reset
			dataa     => add_frame_add_frame_module_frame_parameter_0_vertex_row_wire, --      dataa.wire
			datab     => add_frame_add_frame_module_frame_parameter_0_height_wire,     --      datab.wire
			result    => pipelined_adder1_result_wire,                                 --     result.wire
			user_aclr => pipelined_adder1user_aclrgnd_output_wire,                     --  user_aclr.wire
			ena       => pipelined_adder1enavcc_output_wire                            --        ena.wire
		);

	pipelined_adder1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder1user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder1enavcc_output_wire  -- output.wire
		);

	pipelined_adder2 : component alt_dspbuilder_pipelined_adder_GNWEIMU3MK
		generic map (
			width    => 16,
			pipeline => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => pipelined_adder3_result_wire,             --      dataa.wire
			datab     => constant1_output_wire,                    --      datab.wire
			result    => pipelined_adder2_result_wire,             --     result.wire
			user_aclr => pipelined_adder2user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder2enavcc_output_wire        --        ena.wire
		);

	pipelined_adder2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder2user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder2enavcc_output_wire  -- output.wire
		);

	writedata_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => writedata,               --  input.wire
			output => writedata_0_output_wire  -- output.wire
		);

	constant6 : component alt_dspbuilder_constant_GNWFCSDEFM
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000000000000001",
			width      => 16
		)
		port map (
			output => constant6_output_wire  -- output.wire
		);

	constant7 : component alt_dspbuilder_constant_GNLMV7GZFA
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "111111111111111111111111",
			width      => 24
		)
		port map (
			output => constant7_output_wire  -- output.wire
		);

	addr_0 : component alt_dspbuilder_port_GNS2GDLO5E
		port map (
			input  => addr,               --  input.wire
			output => addr_0_output_wire  -- output.wire
		);

	constant4 : component alt_dspbuilder_constant_GNZEH3JAKA
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000001111",
			width      => 24
		)
		port map (
			output => constant4_output_wire  -- output.wire
		);

	constant5 : component alt_dspbuilder_constant_GNNKZSYI73
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000000",
			width      => 24
		)
		port map (
			output => constant5_output_wire  -- output.wire
		);

	constant8 : component alt_dspbuilder_constant_GNWFCSDEFM
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000000000000001",
			width      => 16
		)
		port map (
			output => constant8_output_wire  -- output.wire
		);

	constant9 : component alt_dspbuilder_constant_GNGITJD4MB
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000011111111",
			width      => 24
		)
		port map (
			output => constant9_output_wire  -- output.wire
		);

	logical_bit_operator7 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator7_result_wire, -- result.wire
			data0  => cast19_output_wire,                --  data0.wire
			data1  => if_statement_true_wire             --  data1.wire
		);

	logical_bit_operator6 : component alt_dspbuilder_logical_bit_op_GN5A3KLAEC
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 3
		)
		port map (
			result => logical_bit_operator6_result_wire, -- result.wire
			data0  => cast18_output_wire,                --  data0.wire
			data1  => if_statement2_true_wire,           --  data1.wire
			data2  => valid_0_output_wire                --  data2.wire
		);

	logical_bit_operator5 : component alt_dspbuilder_logical_bit_op_GNKUBZL4TE
		generic map (
			LogicalOp     => "AltNOT",
			number_inputs => 1
		)
		port map (
			result => logical_bit_operator5_result_wire, -- result.wire
			data0  => cast17_output_wire                 --  data0.wire
		);

	logical_bit_operator4 : component alt_dspbuilder_logical_bit_op_GNUQ2R64DV
		generic map (
			LogicalOp     => "AltOR",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator4_result_wire, -- result.wire
			data0  => if_statement4_true_wire,           --  data0.wire
			data1  => if_statement3_true_wire            --  data1.wire
		);

	constant10 : component alt_dspbuilder_constant_GNNTMI25OE
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000001111111100000000",
			width      => 24
		)
		port map (
			output => constant10_output_wire  -- output.wire
		);

	constant3 : component alt_dspbuilder_constant_GNNKZSYI73
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000000",
			width      => 24
		)
		port map (
			output => constant3_output_wire  -- output.wire
		);

	constant11 : component alt_dspbuilder_constant_GNIJTURCWG
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "111111110000000000000000",
			width      => 24
		)
		port map (
			output => constant11_output_wire  -- output.wire
		);

	if_statement : component alt_dspbuilder_if_statement_GNHRNNRV37
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "(((a>b) or (a=b)) and ((a<c) or (a=c)) and (d=e)) or ((d>e) and (d<f) and (a=b)) or ((d>e) and (d<f) and (a=c)) or (((a>b) or (a=b)) and ((a<c) or (a=c)) and (d=f))",
			number_inputs   => 6,
			width           => 16
		)
		port map (
			true => if_statement_true_wire,                                       -- true.wire
			a    => counter_q_wire,                                               --    a.wire
			b    => add_frame_add_frame_module_frame_parameter_0_vertex_col_wire, --    b.wire
			c    => pipelined_adder_result_wire,                                  --    c.wire
			d    => counter1_q_wire,                                              --    d.wire
			e    => add_frame_add_frame_module_frame_parameter_0_vertex_row_wire, --    e.wire
			f    => pipelined_adder1_result_wire                                  --    f.wire
		);

	constant1 : component alt_dspbuilder_constant_GNWFCSDEFM
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000000000000001",
			width      => 16
		)
		port map (
			output => constant1_output_wire  -- output.wire
		);

	add_frame_add_frame_module_frame_parameter_0 : component Add_Frame_GN_Add_Frame_Add_Frame_Module_FRAME_PARAMETER
		port map (
			writedata  => writedata_0_output_wire,                                      --  writedata.wire
			data       => data_in_0_output_wire,                                        --       data.wire
			height     => add_frame_add_frame_module_frame_parameter_0_height_wire,     --     height.wire
			Clock      => clock_0_clock_output_clk,                                     --      Clock.clk
			aclr       => clock_0_clock_output_reset,                                   --           .reset
			write      => write_0_output_wire,                                          --      write.wire
			width      => add_frame_add_frame_module_frame_parameter_0_width_wire,      --      width.wire
			sop        => sop_0_output_wire,                                            --        sop.wire
			enble      => add_frame_add_frame_module_frame_parameter_0_enble_wire,      --      enble.wire
			addr       => addr_0_output_wire,                                           --       addr.wire
			color      => add_frame_add_frame_module_frame_parameter_0_color_wire,      --      color.wire
			vertex_col => add_frame_add_frame_module_frame_parameter_0_vertex_col_wire, -- vertex_col.wire
			vertex_row => add_frame_add_frame_module_frame_parameter_0_vertex_row_wire  -- vertex_row.wire
		);

	add_frame_add_frame_module_ctrl_decoder_0 : component Add_Frame_GN_Add_Frame_Add_Frame_Module_CTRL_DECODER
		port map (
			height => add_frame_add_frame_module_ctrl_decoder_0_height_wire, -- height.wire
			width  => add_frame_add_frame_module_ctrl_decoder_0_width_wire,  --  width.wire
			sop    => sop_0_output_wire,                                     --    sop.wire
			Clock  => clock_0_clock_output_clk,                              --  Clock.clk
			aclr   => clock_0_clock_output_reset,                            --       .reset
			data   => multiplexer1_result_wire,                              --   data.wire
			valid  => valid_0_output_wire                                    --  valid.wire
		);

	single_pulse : component alt_dspbuilder_single_pulse_GN2XGKTRR3
		generic map (
			delay         => 1,
			signal_type   => "Step Down",
			impulse_width => 1
		)
		port map (
			clock  => clock_0_clock_output_clk,        -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,      --           .reset
			result => single_pulse_result_wire,        --     result.wire
			sclr   => single_pulsesclrgnd_output_wire, --       sclr.wire
			ena    => single_pulseenavcc_output_wire   --        ena.wire
		);

	single_pulsesclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => single_pulsesclrgnd_output_wire  -- output.wire
		);

	single_pulseenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => single_pulseenavcc_output_wire  -- output.wire
		);

	write_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => write,               --  input.wire
			output => write_0_output_wire  -- output.wire
		);

	logical_bit_operator3 : component alt_dspbuilder_logical_bit_op_GNKUBZL4TE
		generic map (
			LogicalOp     => "AltNOT",
			number_inputs => 1
		)
		port map (
			result => logical_bit_operator3_result_wire, -- result.wire
			data0  => cast16_output_wire                 --  data0.wire
		);

	logical_bit_operator2 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator2_result_wire, -- result.wire
			data0  => eop_0_output_wire,                 --  data0.wire
			data1  => cast14_output_wire                 --  data1.wire
		);

	eop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => eop,               --  input.wire
			output => eop_0_output_wire  -- output.wire
		);

	logical_bit_operator1 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator1_result_wire, -- result.wire
			data0  => cast13_output_wire,                --  data0.wire
			data1  => valid_0_output_wire                --  data1.wire
		);

	logical_bit_operator : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator_result_wire, -- result.wire
			data0  => if_statement1_true_wire,          --  data0.wire
			data1  => sop_0_output_wire                 --  data1.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GNTWZRTG4I
		generic map (
			width    => 16,
			pipeline => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,                                     -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                                   --           .reset
			dataa     => add_frame_add_frame_module_frame_parameter_0_vertex_col_wire, --      dataa.wire
			datab     => add_frame_add_frame_module_frame_parameter_0_width_wire,      --      datab.wire
			result    => pipelined_adder_result_wire,                                  --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire,                      --  user_aclr.wire
			ena       => pipelined_adderenavcc_output_wire                             --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adderenavcc_output_wire  -- output.wire
		);

	if_statement4 : component alt_dspbuilder_if_statement_GNUCFELPE2
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "(a=b)",
			number_inputs   => 2,
			width           => 16
		)
		port map (
			true => if_statement4_true_wire,      -- true.wire
			a    => pipelined_adder4_result_wire, --    a.wire
			b    => counter1_q_wire               --    b.wire
		);

	if_statement3 : component alt_dspbuilder_if_statement_GNUCFELPE2
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "(a=b)",
			number_inputs   => 2,
			width           => 16
		)
		port map (
			true => if_statement3_true_wire,      -- true.wire
			a    => pipelined_adder3_result_wire, --    a.wire
			b    => counter_q_wire                --    b.wire
		);

	counter : component alt_dspbuilder_counter_GNCXSYJEM5
		generic map (
			use_usr_aclr => "false",
			use_ena      => "false",
			use_cin      => "false",
			use_sset     => "false",
			ndirection   => 1,
			svalue       => "1",
			use_sload    => "false",
			use_sclr     => "true",
			use_cout     => "false",
			modulus      => -1,
			use_cnt_ena  => "true",
			width        => 16,
			use_aset     => "false",
			use_aload    => "false",
			avalue       => "0"
		)
		port map (
			clock   => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr    => clock_0_clock_output_reset,        --           .reset
			cnt_ena => logical_bit_operator1_result_wire, --    cnt_ena.wire
			sclr    => logical_bit_operator4_result_wire, --       sclr.wire
			q       => counter_q_wire,                    --          q.wire
			cout    => open                               --       cout.wire
		);

	if_statement2 : component alt_dspbuilder_if_statement_GNUCFELPE2
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "(a=b)",
			number_inputs   => 2,
			width           => 16
		)
		port map (
			true => if_statement2_true_wire,      -- true.wire
			a    => pipelined_adder2_result_wire, --    a.wire
			b    => counter_q_wire                --    b.wire
		);

	if_statement1 : component alt_dspbuilder_if_statement_GN7VA7SRUP
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "(a=b) and (a /= c)",
			number_inputs   => 3,
			width           => 24
		)
		port map (
			true => if_statement1_true_wire, -- true.wire
			a    => data_in_0_output_wire,   --    a.wire
			b    => constant3_output_wire,   --    b.wire
			c    => constant4_output_wire    --    c.wire
		);

	frame_control : component FrameControl
		port map (
			clock    => clock_0_clock_output_clk,          --    clock.clk
			reset    => single_pulse_result_wire,          --    reset.wire
			ctrl_in  => logical_bit_operator3_result_wire, --  ctrl_in.wire
			data_in  => cast11_output_wire,                --  data_in.wire
			frame_in => logical_bit_operator7_result_wire, -- frame_in.wire
			state    => frame_control_state_wire           --    state.wire
		);

	delay3 : component alt_dspbuilder_delay_GNHYCSAEGT
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "0",
			width      => 1
		)
		port map (
			input  => cast12_output_wire,         --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay3_output_wire,         --     output.wire
			sclr   => delay3sclrgnd_output_wire,  --       sclr.wire
			ena    => delay3enavcc_output_wire    --        ena.wire
		);

	delay3sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay3sclrgnd_output_wire  -- output.wire
		);

	delay3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay3enavcc_output_wire  -- output.wire
		);

	sop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sop,               --  input.wire
			output => sop_0_output_wire  -- output.wire
		);

	multiplexer1 : component alt_dspbuilder_multiplexer_GNRF25WCVA
		generic map (
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 1,
			width                  => 24,
			pipeline               => 0,
			number_inputs          => 3
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast20_output_wire,                   --        sel.wire
			result    => multiplexer1_result_wire,             --     result.wire
			ena       => multiplexer1enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer1user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => data_in_0_output_wire,                --        in0.wire
			in1       => data_in_0_output_wire,                --        in1.wire
			in2       => multiplexer2_result_wire              --        in2.wire
		);

	multiplexer1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer1user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer1enavcc_output_wire  -- output.wire
		);

	delay1 : component alt_dspbuilder_delay_GNUECIBFDH
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "0",
			width      => 1
		)
		port map (
			input  => delay3_output_wire,         --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay1_output_wire,         --     output.wire
			sclr   => cast9_output_wire,          --       sclr.wire
			ena    => cast10_output_wire          --        ena.wire
		);

	multiplexer2 : component alt_dspbuilder_multiplexer_GNHHROOGAI
		generic map (
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0,
			width                  => 24,
			pipeline               => 0,
			number_inputs          => 5
		)
		port map (
			clock     => clock_0_clock_output_clk,                                -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                              --           .reset
			sel       => add_frame_add_frame_module_frame_parameter_0_color_wire, --        sel.wire
			result    => multiplexer2_result_wire,                                --     result.wire
			ena       => multiplexer2enavcc_output_wire,                          --        ena.wire
			user_aclr => multiplexer2user_aclrgnd_output_wire,                    --  user_aclr.wire
			in0       => constant5_output_wire,                                   --        in0.wire
			in1       => constant7_output_wire,                                   --        in1.wire
			in2       => constant9_output_wire,                                   --        in2.wire
			in3       => constant10_output_wire,                                  --        in3.wire
			in4       => constant11_output_wire                                   --        in4.wire
		);

	multiplexer2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer2user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer2enavcc_output_wire  -- output.wire
		);

	delay2 : component alt_dspbuilder_delay_GNHYCSAEGT
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "0",
			width      => 1
		)
		port map (
			input  => cast15_output_wire,         --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay2_output_wire,         --     output.wire
			sclr   => delay2sclrgnd_output_wire,  --       sclr.wire
			ena    => delay2enavcc_output_wire    --        ena.wire
		);

	delay2sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay2sclrgnd_output_wire  -- output.wire
		);

	delay2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay2enavcc_output_wire  -- output.wire
		);

	data_out_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => multiplexer1_result_wire, --  input.wire
			output => data_out                  -- output.wire
		);

	data_in_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => data_in,               --  input.wire
			output => data_in_0_output_wire  -- output.wire
		);

	counter1 : component alt_dspbuilder_counter_GNCXSYJEM5
		generic map (
			use_usr_aclr => "false",
			use_ena      => "false",
			use_cin      => "false",
			use_sset     => "false",
			ndirection   => 1,
			svalue       => "1",
			use_sload    => "false",
			use_sclr     => "true",
			use_cout     => "false",
			modulus      => -1,
			use_cnt_ena  => "true",
			width        => 16,
			use_aset     => "false",
			use_aload    => "false",
			avalue       => "0"
		)
		port map (
			clock   => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr    => clock_0_clock_output_reset,        --           .reset
			cnt_ena => logical_bit_operator6_result_wire, --    cnt_ena.wire
			sclr    => logical_bit_operator5_result_wire, --       sclr.wire
			q       => counter1_q_wire,                   --          q.wire
			cout    => open                               --       cout.wire
		);

	cast9 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay2_output_wire, --  input.wire
			output => cast9_output_wire   -- output.wire
		);

	cast10 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay3_output_wire, --  input.wire
			output => cast10_output_wire  -- output.wire
		);

	cast11 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire, --  input.wire
			output => cast11_output_wire  -- output.wire
		);

	cast12 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator_result_wire, --  input.wire
			output => cast12_output_wire                -- output.wire
		);

	cast13 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire, --  input.wire
			output => cast13_output_wire  -- output.wire
		);

	cast14 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire, --  input.wire
			output => cast14_output_wire  -- output.wire
		);

	cast15 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bit_operator2_result_wire, --  input.wire
			output => cast15_output_wire                 -- output.wire
		);

	cast16 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire, --  input.wire
			output => cast16_output_wire  -- output.wire
		);

	cast17 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire, --  input.wire
			output => cast17_output_wire  -- output.wire
		);

	cast18 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay1_output_wire, --  input.wire
			output => cast18_output_wire  -- output.wire
		);

	cast19 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => add_frame_add_frame_module_frame_parameter_0_enble_wire, --  input.wire
			output => cast19_output_wire                                       -- output.wire
		);

	cast20 : component alt_dspbuilder_cast_GNLWRZWTQF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => frame_control_state_wire, --  input.wire
			output => cast20_output_wire        -- output.wire
		);

end architecture rtl; -- of Add_Frame_GN_Add_Frame_Add_Frame_Module
