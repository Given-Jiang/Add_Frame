-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Full Version
-- Created on Sun Feb 22 16:00:27 2015

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FrameControl IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        ctrl_in : IN STD_LOGIC := '0';
        data_in : IN STD_LOGIC := '0';
        frame_in : IN STD_LOGIC := '0';
        state : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
    );
END FrameControl;

ARCHITECTURE BEHAVIOR OF FrameControl IS
    TYPE type_fstate IS (IDLE,DATA,FRAME,CTRL);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,ctrl_in,data_in,frame_in)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= IDLE;
            state <= "000";
        ELSE
            state <= "000";
            CASE fstate IS
                WHEN IDLE =>
                    IF ((ctrl_in = '1')) THEN
                        reg_fstate <= CTRL;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= IDLE;
                    END IF;

                    state <= "000";
                WHEN DATA =>
                    IF (((ctrl_in = '0') AND (frame_in = '1'))) THEN
                        reg_fstate <= FRAME;
                    ELSIF (((ctrl_in = '1') AND (frame_in = '0'))) THEN
                        reg_fstate <= CTRL;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= DATA;
                    END IF;

                    state <= "010";
                WHEN FRAME =>
                    IF ((((ctrl_in = '1') AND (data_in = '0')) AND (frame_in = '0'))) THEN
                        reg_fstate <= CTRL;
                    ELSIF ((((ctrl_in = '0') AND (data_in = '1')) AND (frame_in = '0'))) THEN
                        reg_fstate <= DATA;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= FRAME;
                    END IF;

                    state <= "100";
                WHEN CTRL =>
                    IF (((data_in = '0') AND (frame_in = '1'))) THEN
                        reg_fstate <= FRAME;
                    ELSIF (((data_in = '1') AND (frame_in = '0'))) THEN
                        reg_fstate <= DATA;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= CTRL;
                    END IF;

                    state <= "001";
                WHEN OTHERS => 
                    state <= "XXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
